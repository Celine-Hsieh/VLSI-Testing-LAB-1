
module c499 ( xid0, xid1, xid2, xid3, xid4, xid5, xid6, xid7, xid8, xid9, 
        xid10, xid11, xid12, xid13, xid14, xid15, xid16, xid17, xid18, xid19, 
        xid20, xid21, xid22, xid23, xid24, xid25, xid26, xid27, xid28, xid29, 
        xid30, xid31, xic0, xic1, xic2, xic3, xic4, xic5, xic6, xic7, xr, xod0, 
        xod1, xod2, xod3, xod4, xod5, xod6, xod7, xod8, xod9, xod10, xod11, 
        xod12, xod13, xod14, xod15, xod16, xod17, xod18, xod19, xod20, xod21, 
        xod22, xod23, xod24, xod25, xod26, xod27, xod28, xod29, xod30, xod31
 );
  input xid0, xid1, xid2, xid3, xid4, xid5, xid6, xid7, xid8, xid9, xid10,
         xid11, xid12, xid13, xid14, xid15, xid16, xid17, xid18, xid19, xid20,
         xid21, xid22, xid23, xid24, xid25, xid26, xid27, xid28, xid29, xid30,
         xid31, xic0, xic1, xic2, xic3, xic4, xic5, xic6, xic7, xr;
  output xod0, xod1, xod2, xod3, xod4, xod5, xod6, xod7, xod8, xod9, xod10,
         xod11, xod12, xod13, xod14, xod15, xod16, xod17, xod18, xod19, xod20,
         xod21, xod22, xod23, xod24, xod25, xod26, xod27, xod28, xod29, xod30,
         xod31;
  wire   n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281;

  XNOR2X1 U178 ( .A(xid9), .B(n146), .Y(xod9) );
  NAND2X1 U179 ( .A(n147), .B(n148), .Y(n146) );
  XNOR2X1 U180 ( .A(xid8), .B(n149), .Y(xod8) );
  NAND2X1 U181 ( .A(n147), .B(n150), .Y(n149) );
  XNOR2X1 U182 ( .A(xid7), .B(n151), .Y(xod7) );
  NAND2X1 U183 ( .A(n152), .B(n153), .Y(n151) );
  XNOR2X1 U184 ( .A(xid6), .B(n154), .Y(xod6) );
  NAND2X1 U185 ( .A(n152), .B(n155), .Y(n154) );
  XNOR2X1 U186 ( .A(xid5), .B(n156), .Y(xod5) );
  NAND2X1 U187 ( .A(n152), .B(n148), .Y(n156) );
  XNOR2X1 U188 ( .A(xid4), .B(n157), .Y(xod4) );
  NAND2X1 U189 ( .A(n152), .B(n150), .Y(n157) );
  AND4X1 U190 ( .A(n158), .B(n159), .C(n160), .D(n161), .Y(n152) );
  XNOR2X1 U191 ( .A(xid31), .B(n162), .Y(xod31) );
  NAND2X1 U192 ( .A(n163), .B(n164), .Y(n162) );
  XNOR2X1 U193 ( .A(xid30), .B(n165), .Y(xod30) );
  NAND2X1 U194 ( .A(n163), .B(n166), .Y(n165) );
  XNOR2X1 U195 ( .A(xid3), .B(n167), .Y(xod3) );
  NAND2X1 U196 ( .A(n168), .B(n153), .Y(n167) );
  XNOR2X1 U197 ( .A(xid29), .B(n169), .Y(xod29) );
  NAND2X1 U198 ( .A(n163), .B(n170), .Y(n169) );
  XNOR2X1 U199 ( .A(xid28), .B(n171), .Y(xod28) );
  NAND2X1 U200 ( .A(n163), .B(n172), .Y(n171) );
  AND4X1 U201 ( .A(n148), .B(n173), .C(n153), .D(n174), .Y(n163) );
  NOR2X1 U202 ( .A(n155), .B(n150), .Y(n174) );
  XNOR2X1 U203 ( .A(xid27), .B(n175), .Y(xod27) );
  NAND2X1 U204 ( .A(n176), .B(n164), .Y(n175) );
  XNOR2X1 U205 ( .A(xid26), .B(n177), .Y(xod26) );
  NAND2X1 U206 ( .A(n176), .B(n166), .Y(n177) );
  XNOR2X1 U207 ( .A(xid25), .B(n178), .Y(xod25) );
  NAND2X1 U208 ( .A(n176), .B(n170), .Y(n178) );
  XNOR2X1 U209 ( .A(xid24), .B(n179), .Y(xod24) );
  NAND2X1 U210 ( .A(n176), .B(n172), .Y(n179) );
  AND4X1 U211 ( .A(n180), .B(n181), .C(n182), .D(n173), .Y(n176) );
  XNOR2X1 U212 ( .A(xid23), .B(n183), .Y(xod23) );
  NAND2X1 U213 ( .A(n184), .B(n164), .Y(n183) );
  XNOR2X1 U214 ( .A(xid22), .B(n185), .Y(xod22) );
  NAND2X1 U215 ( .A(n184), .B(n166), .Y(n185) );
  XNOR2X1 U216 ( .A(xid21), .B(n186), .Y(xod21) );
  NAND2X1 U217 ( .A(n184), .B(n170), .Y(n186) );
  XNOR2X1 U218 ( .A(xid20), .B(n187), .Y(xod20) );
  NAND2X1 U219 ( .A(n184), .B(n172), .Y(n187) );
  AND4X1 U220 ( .A(n188), .B(n189), .C(n190), .D(n173), .Y(n184) );
  XNOR2X1 U221 ( .A(xid2), .B(n191), .Y(xod2) );
  NAND2X1 U222 ( .A(n168), .B(n155), .Y(n191) );
  XNOR2X1 U223 ( .A(xid19), .B(n192), .Y(xod19) );
  NAND2X1 U224 ( .A(n193), .B(n164), .Y(n192) );
  XNOR2X1 U225 ( .A(xid18), .B(n194), .Y(xod18) );
  NAND2X1 U226 ( .A(n193), .B(n166), .Y(n194) );
  XNOR2X1 U227 ( .A(xid17), .B(n195), .Y(xod17) );
  NAND2X1 U228 ( .A(n193), .B(n170), .Y(n195) );
  XNOR2X1 U229 ( .A(xid16), .B(n196), .Y(xod16) );
  NAND2X1 U230 ( .A(n193), .B(n172), .Y(n196) );
  AND4X1 U231 ( .A(n155), .B(n173), .C(n150), .D(n197), .Y(n193) );
  NOR2X1 U232 ( .A(n148), .B(n153), .Y(n197) );
  OAI33X1 U233 ( .A0(n170), .A1(n159), .A2(n166), .B0(n164), .B1(n198), .B2(
        n172), .Y(n173) );
  AND2X1 U234 ( .A(n172), .B(n164), .Y(n159) );
  XNOR2X1 U235 ( .A(xid15), .B(n199), .Y(xod15) );
  NAND2X1 U236 ( .A(n200), .B(n153), .Y(n199) );
  XNOR2X1 U237 ( .A(xid14), .B(n201), .Y(xod14) );
  NAND2X1 U238 ( .A(n200), .B(n155), .Y(n201) );
  XNOR2X1 U239 ( .A(xid13), .B(n202), .Y(xod13) );
  NAND2X1 U240 ( .A(n200), .B(n148), .Y(n202) );
  XNOR2X1 U241 ( .A(xid12), .B(n203), .Y(xod12) );
  NAND2X1 U242 ( .A(n200), .B(n150), .Y(n203) );
  AND4X1 U243 ( .A(n164), .B(n161), .C(n170), .D(n204), .Y(n200) );
  NOR2X1 U244 ( .A(n172), .B(n166), .Y(n204) );
  XNOR2X1 U245 ( .A(xid11), .B(n205), .Y(xod11) );
  NAND2X1 U246 ( .A(n147), .B(n153), .Y(n205) );
  XNOR2X1 U247 ( .A(xid10), .B(n206), .Y(xod10) );
  NAND2X1 U248 ( .A(n147), .B(n155), .Y(n206) );
  NOR4BBX1 U249 ( .AN(n161), .BN(n198), .C(n164), .D(n172), .Y(n147) );
  NOR2X1 U250 ( .A(n160), .B(n158), .Y(n198) );
  CLKINVX1 U251 ( .A(n170), .Y(n158) );
  CLKINVX1 U252 ( .A(n166), .Y(n160) );
  XNOR2X1 U253 ( .A(xid1), .B(n207), .Y(xod1) );
  NAND2X1 U254 ( .A(n168), .B(n148), .Y(n207) );
  XNOR2X1 U255 ( .A(xid0), .B(n208), .Y(xod0) );
  NAND2X1 U256 ( .A(n168), .B(n150), .Y(n208) );
  AND4X1 U257 ( .A(n172), .B(n161), .C(n166), .D(n209), .Y(n168) );
  NOR2X1 U258 ( .A(n164), .B(n170), .Y(n209) );
  XNOR2X1 U259 ( .A(n210), .B(n211), .Y(n170) );
  XOR2X1 U260 ( .A(n212), .B(n213), .Y(n211) );
  XOR2X1 U261 ( .A(xid21), .B(xid17), .Y(n213) );
  XOR2X1 U262 ( .A(xid29), .B(xid25), .Y(n212) );
  XOR2X1 U263 ( .A(n214), .B(n215), .Y(n210) );
  XOR2X1 U264 ( .A(n216), .B(n217), .Y(n214) );
  NAND2X1 U265 ( .A(xic5), .B(xr), .Y(n216) );
  XNOR2X1 U266 ( .A(n218), .B(n219), .Y(n164) );
  XOR2X1 U267 ( .A(n220), .B(n221), .Y(n219) );
  XOR2X1 U268 ( .A(xid23), .B(xid19), .Y(n221) );
  XOR2X1 U269 ( .A(xid31), .B(xid27), .Y(n220) );
  XOR2X1 U270 ( .A(n222), .B(n217), .Y(n218) );
  XNOR2X1 U271 ( .A(n223), .B(n224), .Y(n217) );
  XOR2X1 U272 ( .A(xid15), .B(xid14), .Y(n224) );
  XNOR2X1 U273 ( .A(xid12), .B(xid13), .Y(n223) );
  XOR2X1 U274 ( .A(n225), .B(n226), .Y(n222) );
  NAND2X1 U275 ( .A(xic7), .B(xr), .Y(n225) );
  XNOR2X1 U276 ( .A(n227), .B(n228), .Y(n166) );
  XOR2X1 U277 ( .A(n229), .B(n230), .Y(n228) );
  XOR2X1 U278 ( .A(xid22), .B(xid18), .Y(n230) );
  XOR2X1 U279 ( .A(xid30), .B(xid26), .Y(n229) );
  XOR2X1 U280 ( .A(n231), .B(n215), .Y(n227) );
  XNOR2X1 U281 ( .A(n232), .B(n233), .Y(n215) );
  XOR2X1 U282 ( .A(xid9), .B(xid8), .Y(n233) );
  XNOR2X1 U283 ( .A(xid10), .B(xid11), .Y(n232) );
  XOR2X1 U284 ( .A(n234), .B(n235), .Y(n231) );
  NAND2X1 U285 ( .A(xic6), .B(xr), .Y(n234) );
  OAI33X1 U286 ( .A0(n155), .A1(n189), .A2(n148), .B0(n150), .B1(n181), .B2(
        n153), .Y(n161) );
  NOR2X1 U287 ( .A(n190), .B(n188), .Y(n181) );
  CLKINVX1 U288 ( .A(n155), .Y(n188) );
  CLKINVX1 U289 ( .A(n148), .Y(n190) );
  XNOR2X1 U290 ( .A(n236), .B(n237), .Y(n148) );
  XOR2X1 U291 ( .A(n238), .B(n239), .Y(n237) );
  XOR2X1 U292 ( .A(xid13), .B(xid1), .Y(n239) );
  XOR2X1 U293 ( .A(xid9), .B(xid5), .Y(n238) );
  XOR2X1 U294 ( .A(n240), .B(n241), .Y(n236) );
  XOR2X1 U295 ( .A(n242), .B(n243), .Y(n240) );
  NAND2X1 U296 ( .A(xic1), .B(xr), .Y(n242) );
  NOR2X1 U297 ( .A(n182), .B(n180), .Y(n189) );
  CLKINVX1 U298 ( .A(n150), .Y(n180) );
  XNOR2X1 U299 ( .A(n244), .B(n245), .Y(n150) );
  XOR2X1 U300 ( .A(n246), .B(n247), .Y(n245) );
  XOR2X1 U301 ( .A(xid12), .B(xid0), .Y(n247) );
  XOR2X1 U302 ( .A(xid8), .B(xid4), .Y(n246) );
  XOR2X1 U303 ( .A(n248), .B(n249), .Y(n244) );
  XOR2X1 U304 ( .A(n250), .B(n251), .Y(n248) );
  NAND2X1 U305 ( .A(xic0), .B(xr), .Y(n250) );
  CLKINVX1 U306 ( .A(n153), .Y(n182) );
  XNOR2X1 U307 ( .A(n252), .B(n253), .Y(n153) );
  XOR2X1 U308 ( .A(n254), .B(n255), .Y(n253) );
  XOR2X1 U309 ( .A(xid15), .B(xid11), .Y(n255) );
  XOR2X1 U310 ( .A(xid7), .B(xid3), .Y(n254) );
  XOR2X1 U311 ( .A(n256), .B(n249), .Y(n252) );
  XNOR2X1 U312 ( .A(n257), .B(n258), .Y(n249) );
  XOR2X1 U313 ( .A(xid23), .B(xid22), .Y(n258) );
  XNOR2X1 U314 ( .A(xid20), .B(xid21), .Y(n257) );
  XOR2X1 U315 ( .A(n259), .B(n241), .Y(n256) );
  XNOR2X1 U316 ( .A(n260), .B(n261), .Y(n241) );
  XOR2X1 U317 ( .A(xid31), .B(xid30), .Y(n261) );
  XNOR2X1 U318 ( .A(xid28), .B(xid29), .Y(n260) );
  NAND2X1 U319 ( .A(xic3), .B(xr), .Y(n259) );
  XNOR2X1 U320 ( .A(n262), .B(n263), .Y(n155) );
  XOR2X1 U321 ( .A(n264), .B(n265), .Y(n263) );
  XOR2X1 U322 ( .A(xid14), .B(xid10), .Y(n265) );
  XOR2X1 U323 ( .A(xid6), .B(xid2), .Y(n264) );
  XOR2X1 U324 ( .A(n266), .B(n251), .Y(n262) );
  XNOR2X1 U325 ( .A(n267), .B(n268), .Y(n251) );
  XOR2X1 U326 ( .A(xid19), .B(xid18), .Y(n268) );
  XNOR2X1 U327 ( .A(xid16), .B(xid17), .Y(n267) );
  XOR2X1 U328 ( .A(n269), .B(n243), .Y(n266) );
  XNOR2X1 U329 ( .A(n270), .B(n271), .Y(n243) );
  XOR2X1 U330 ( .A(xid27), .B(xid26), .Y(n271) );
  XNOR2X1 U331 ( .A(xid24), .B(xid25), .Y(n270) );
  NAND2X1 U332 ( .A(xr), .B(xic2), .Y(n269) );
  XNOR2X1 U333 ( .A(n272), .B(n273), .Y(n172) );
  XOR2X1 U334 ( .A(n274), .B(n275), .Y(n273) );
  XOR2X1 U335 ( .A(xid20), .B(xid16), .Y(n275) );
  XOR2X1 U336 ( .A(xid28), .B(xid24), .Y(n274) );
  XOR2X1 U337 ( .A(n276), .B(n226), .Y(n272) );
  XNOR2X1 U338 ( .A(n277), .B(n278), .Y(n226) );
  XOR2X1 U339 ( .A(xid7), .B(xid6), .Y(n278) );
  XNOR2X1 U340 ( .A(xid4), .B(xid5), .Y(n277) );
  XOR2X1 U341 ( .A(n279), .B(n235), .Y(n276) );
  XNOR2X1 U342 ( .A(n280), .B(n281), .Y(n235) );
  XOR2X1 U343 ( .A(xid3), .B(xid2), .Y(n281) );
  XNOR2X1 U344 ( .A(xid0), .B(xid1), .Y(n280) );
  NAND2X1 U345 ( .A(xic4), .B(xr), .Y(n279) );
endmodule

